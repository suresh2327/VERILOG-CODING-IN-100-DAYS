//desgin code for D flip flop
module D_FF(input clk,input d,output reg q);
    always @(posedge clk) begin
        q <= d;
    end
endmodule
